/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  wire load = uio_in[0];
  reg [7:0] value;
  assign uo_out = ena ? value : 8'bzzzzzzzz;

  always @(posedge clk or negedge rst_n) begin
      // asynchronous reset
      if (rst_n == 1'b0) begin
        value <= 8'b00000000;
      // synchronous load
      end else if (load == 1'b1) begin
          value <= ui_in;
      // increment
      end else begin
          value <= value + 1'b1;
      end
  end

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, uio_in [7:1], 1'b0};

endmodule
